// megafunction wizard: %RAM initializer%
// GENERATION: STANDARD
// VERSION: WM1.0
// MODULE: ALTMEM_INIT 

// ============================================================
// File Name: memory.v
// Megafunction Name(s):
// 			ALTMEM_INIT
//
// Simulation Library Files(s):
// 			
// ============================================================
// ************************************************************
// THIS IS A WIZARD-GENERATED FILE. DO NOT EDIT THIS FILE!
//
// 16.0.0 Build 211 04/27/2016 SJ Lite Edition
// ************************************************************


//Copyright (C) 1991-2016 Altera Corporation. All rights reserved.
//Your use of Altera Corporation's design tools, logic functions 
//and other software and tools, and its AMPP partner logic 
//functions, and any output files from any of the foregoing 
//(including device programming or simulation files), and any 
//associated documentation or information are expressly subject 
//to the terms and conditions of the Altera Program License 
//Subscription Agreement, the Altera Quartus Prime License Agreement,
//the Altera MegaCore Function License Agreement, or other 
//applicable license agreement, including, without limitation, 
//that your use is for the sole purpose of programming logic 
//devices manufactured by Altera and sold by Altera or its 
//authorized distributors.  Please refer to the applicable 
//agreement for further details.


// synopsys translate_off
`timescale 1 ps / 1 ps
// synopsys translate_on
module memory (
	clock,
	init,
	dataout,
	init_busy,
	ram_address,
	ram_wren);

	input	  clock;
	input	  init;
	output	[31:0]  dataout;
	output	  init_busy;
	output	[15:0]  ram_address;
	output	  ram_wren;

	wire [31:0] sub_wire0;
	wire  sub_wire1;
	wire [15:0] sub_wire2;
	wire  sub_wire3;
	wire [31:0] dataout = sub_wire0[31:0];
	wire  init_busy = sub_wire1;
	wire [15:0] ram_address = sub_wire2[15:0];
	wire  ram_wren = sub_wire3;

	altmem_init	ALTMEM_INIT_component (
				.clock (clock),
				.init (init),
				.dataout (sub_wire0),
				.init_busy (sub_wire1),
				.ram_address (sub_wire2),
				.ram_wren (sub_wire3),
				.clken (1'b1),
				.datain ({32{1'b0}}),
				.rom_address (),
				.rom_data_ready (1'b0),
				.rom_rden ());
	defparam
		ALTMEM_INIT_component.init_file = "teste1binario8.input",
		ALTMEM_INIT_component.init_to_zero = "NO",
		ALTMEM_INIT_component.intended_device_family = "Cyclone IV E",
		ALTMEM_INIT_component.lpm_hint = "UNUSED",
		ALTMEM_INIT_component.lpm_type = "altmem_init",
		ALTMEM_INIT_component.numwords = 65536,
		ALTMEM_INIT_component.port_rom_data_ready = "PORT_UNUSED",
		ALTMEM_INIT_component.rom_read_latency = 1,
		ALTMEM_INIT_component.width = 32,
		ALTMEM_INIT_component.widthad = 16;


endmodule

// ============================================================
// CNX file retrieval info
// ============================================================
// Retrieval info: LIBRARY: altera_mf altera_mf.altera_mf_components.all
// Retrieval info: PRIVATE: INTENDED_DEVICE_FAMILY STRING "Cyclone IV E"
// Retrieval info: CONSTANT: INIT_FILE STRING "teste1binario8.input"
// Retrieval info: CONSTANT: INIT_TO_ZERO STRING "NO"
// Retrieval info: CONSTANT: INTENDED_DEVICE_FAMILY STRING "Cyclone IV E"
// Retrieval info: CONSTANT: LPM_HINT STRING "UNUSED"
// Retrieval info: CONSTANT: LPM_TYPE STRING "altmem_init"
// Retrieval info: CONSTANT: NUMWORDS NUMERIC "65536"
// Retrieval info: CONSTANT: PORT_ROM_DATA_READY STRING "PORT_UNUSED"
// Retrieval info: CONSTANT: ROM_READ_LATENCY NUMERIC "1"
// Retrieval info: CONSTANT: WIDTH NUMERIC "32"
// Retrieval info: CONSTANT: WIDTHAD NUMERIC "16"
// Retrieval info: USED_PORT: clock 0 0 0 0 INPUT NODEFVAL "clock"
// Retrieval info: CONNECT: @clock 0 0 0 0 clock 0 0 0 0
// Retrieval info: USED_PORT: dataout 0 0 32 0 OUTPUT NODEFVAL "dataout[31..0]"
// Retrieval info: CONNECT: dataout 0 0 32 0 @dataout 0 0 32 0
// Retrieval info: USED_PORT: init 0 0 0 0 INPUT NODEFVAL "init"
// Retrieval info: CONNECT: @init 0 0 0 0 init 0 0 0 0
// Retrieval info: USED_PORT: init_busy 0 0 0 0 OUTPUT NODEFVAL "init_busy"
// Retrieval info: CONNECT: init_busy 0 0 0 0 @init_busy 0 0 0 0
// Retrieval info: USED_PORT: ram_address 0 0 16 0 OUTPUT NODEFVAL "ram_address[15..0]"
// Retrieval info: CONNECT: ram_address 0 0 16 0 @ram_address 0 0 16 0
// Retrieval info: USED_PORT: ram_wren 0 0 0 0 OUTPUT NODEFVAL "ram_wren"
// Retrieval info: CONNECT: ram_wren 0 0 0 0 @ram_wren 0 0 0 0
// Retrieval info: GEN_FILE: TYPE_NORMAL memory.v TRUE FALSE
// Retrieval info: GEN_FILE: TYPE_NORMAL memory.qip TRUE FALSE
// Retrieval info: GEN_FILE: TYPE_NORMAL memory.bsf FALSE TRUE
// Retrieval info: GEN_FILE: TYPE_NORMAL memory_inst.v FALSE TRUE
// Retrieval info: GEN_FILE: TYPE_NORMAL memory_bb.v FALSE TRUE
// Retrieval info: GEN_FILE: TYPE_NORMAL memory.inc FALSE TRUE
// Retrieval info: GEN_FILE: TYPE_NORMAL memory.cmp FALSE TRUE
