//------------------------------------------------------------------------------
//	Module:		LevelToPulse
//	Desc:		This module provides a 1-cycle output based on a push button
//				raw input source.
//	Params:		This module is not parameterized.
//	Inputs:		See Lab2 document
//	Outputs:	See Lab2 document
//
//	Author:     YOUR NAME GOES HERE
//------------------------------------------------------------------------------
module	LevelToPulse(
			//------------------------------------------------------------------
			//	Clock & Reset Inputs
			//------------------------------------------------------------------
			Clock,
			Reset,
			//------------------------------------------------------------------
			
			//------------------------------------------------------------------
			//	Inputs
			//------------------------------------------------------------------
			Level,
			//------------------------------------------------------------------
			
			//------------------------------------------------------------------
			//	Outputs
			//------------------------------------------------------------------
			Pulse
			//------------------------------------------------------------------
	);
	//--------------------------------------------------------------------------
	//	Clock & Reset Inputs
	//--------------------------------------------------------------------------
	input					Clock;	// System clock
	input					Reset;	// System reset
	//--------------------------------------------------------------------------
	
	//--------------------------------------------------------------------------
	//	Inputs
	//--------------------------------------------------------------------------
	input					Level;
	//--------------------------------------------------------------------------

	//--------------------------------------------------------------------------
	//	Outputs
	//--------------------------------------------------------------------------
	output					Pulse;
	//--------------------------------------------------------------------------

	//--------------------------------------------------------------------------
	//	State Encoding
	//--------------------------------------------------------------------------
	
	localparam ativado =1 'b1,
				desativado = 1'b0;

	reg state,next;
	
	//--------------------------------------------------------------------------
	
	//--------------------------------------------------------------------------
	//	Wire Declarations
	//--------------------------------------------------------------------------
	
	// place wire declarations here	
	
	//--------------------------------------------------------------------------
	
	//--------------------------------------------------------------------------
	//	Logic
	//--------------------------------------------------------------------------
	always @(posedge Clock)
		begin
			state <= desativado;
		end
		
	always @(state or Level or Reset) 
		begin
			case(state)
				desativado:
					begin
						Pulse = 1'b0;
						if(Level and !Reset)
							next = ativado;
						else
							next = desativado;
					end
				ativado: 
					begin 
						Pulse = 1'b1;
						next = desativado;
					end
			endcase
		end
	// Place you *behavioral* Verilog here
	// You may find it useful to use a case statement to describe your FSM.

	//--------------------------------------------------------------------------
endmodule // LevelToPulse