//------------------------------------------------------------------------------
//	Module:		LevelToPulse
//	Desc:		This module provides a 1-cycle output based on a push button
//				raw input source.
//	Params:		This module is not parameterized.
//	Inputs:		See Lab2 document
//	Outputs:	See Lab2 document
//
//	Author:     YOUR NAME GOES HERE
//------------------------------------------------------------------------------
module	LevelToPulse(
			//------------------------------------------------------------------
			//	Clock & Reset Inputs
			//------------------------------------------------------------------
			Clock,
			Reset,
			//------------------------------------------------------------------
			
			//------------------------------------------------------------------
			//	Inputs
			//------------------------------------------------------------------
			Level,
			//------------------------------------------------------------------
			
			//------------------------------------------------------------------
			//	Outputs
			//------------------------------------------------------------------
			Pulse
			//------------------------------------------------------------------
	);
	//--------------------------------------------------------------------------
	//	Clock & Reset Inputs
	//--------------------------------------------------------------------------
	input					Clock;	// System clock
	input					Reset;	// System reset
	//--------------------------------------------------------------------------
	
	//--------------------------------------------------------------------------
	//	Inputs
	//--------------------------------------------------------------------------
	input					Level;
	//--------------------------------------------------------------------------

	//--------------------------------------------------------------------------
	//	Outputs
	//--------------------------------------------------------------------------
	output					Pulse;
	//--------------------------------------------------------------------------

	//--------------------------------------------------------------------------
	//	State Encoding
	//--------------------------------------------------------------------------
	
	// place state encoding here
	
	//--------------------------------------------------------------------------
	
	//--------------------------------------------------------------------------
	//	Wire Declarations
	//--------------------------------------------------------------------------
	
	// place wire declarations here	
	
	//--------------------------------------------------------------------------
	
	//--------------------------------------------------------------------------
	//	Logic
	//--------------------------------------------------------------------------
	
	// Place you *behavioral* Verilog here
	// You may find it useful to use a case statement to describe your FSM.

	//--------------------------------------------------------------------------
endmodule // LevelToPulse